module Cor (x, y, a);
input x, y;

output a;


assign a = x | y;

endmodule
