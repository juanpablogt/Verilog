module modulo1 (s,c,a,b);

input a,b;
output s,c;

assign s = a ^ b;
output  c = a & b;

endmodule

